`timescale 1ns / 1ps

module mux2_1_gates(
    input A,
    input B,
    input SEL,
    output OUT
    );


endmodule
