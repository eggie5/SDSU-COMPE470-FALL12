`timescale 1ns / 1ps

module adder_1_bit(
    input A,
    input B,
    output SUM
    );

	assign SUM = A+B;

endmodule
